intiial begin
	a = 5;
	b = 2;

	a <= b;
	b <= a;
end