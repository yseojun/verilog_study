// a===b, a!==b; -> 1,0,z,x 의 logical equallity 판단
